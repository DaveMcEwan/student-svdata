module test (
    input a /* kommentar till port */ /* a */
    );
endmodule